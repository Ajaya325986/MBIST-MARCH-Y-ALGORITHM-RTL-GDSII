* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : controller1                                  *
* Netlisted  : Tue Nov 26 12:01:54 2024                     *
* PVS Version: 22.20-p031 Thu Nov 17 19:06:38 PST 2022      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(nmos1v) _nmos_12 ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(pmos1v) _pmos_12 pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND3BX1                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND3BX1 Y C B VDD VSS AN
** N=9 EP=6 FDC=8
M0 8 C Y VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=1110 $Y=800 $dt=0
M1 9 B 8 VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=1550 $Y=800 $dt=0
M2 VSS 7 9 VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=2190 $Y=800 $dt=0
M3 7 AN VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3150 $Y=1180 $dt=0
M4 VDD C Y VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=710 $Y=3120 $dt=1
M5 Y B VDD VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=1550 $Y=3120 $dt=1
M6 VDD 7 Y VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=2390 $Y=3120 $dt=1
M7 7 AN VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3350 $Y=3120 $dt=1
.ends NAND3BX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: CLKINVX1                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt CLKINVX1 A Y VDD VSS
** N=4 EP=4 FDC=2
M0 Y A VSS VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=710 $Y=870 $dt=0
M1 Y A VDD VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=710 $Y=2680 $dt=1
.ends CLKINVX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OAI211XL                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OAI211XL A1 B0 A0 Y VDD VSS C0
** N=10 EP=7 FDC=8
M0 VSS A0 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=710 $Y=1140 $dt=0
M1 8 A1 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1550 $Y=1140 $dt=0
M2 9 B0 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2390 $Y=1140 $dt=0
M3 Y C0 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2830 $Y=1140 $dt=0
M4 10 A0 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=820 $Y=3180 $dt=1
M5 Y A1 10 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1260 $Y=3180 $dt=1
M6 VDD B0 Y VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2100 $Y=3180 $dt=1
M7 Y C0 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3150 $Y=3180 $dt=1
.ends OAI211XL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AOI211XL                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AOI211XL A1 B0 A0 Y VDD VSS C0
** N=10 EP=7 FDC=8
M0 8 A0 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=710 $Y=1030 $dt=0
M1 Y A1 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1150 $Y=1030 $dt=0
M2 VSS B0 Y VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1990 $Y=1030 $dt=0
M3 Y C0 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2830 $Y=1030 $dt=0
M4 VDD A0 9 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=710 $Y=3380 $dt=1
M5 9 A1 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1550 $Y=3380 $dt=1
M6 10 B0 9 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2390 $Y=3380 $dt=1
M7 Y C0 10 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2830 $Y=3380 $dt=1
.ends AOI211XL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OAI21XL                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OAI21XL A1 A0 VDD VSS B0 Y
** N=8 EP=6 FDC=6
M0 VSS A0 7 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=890 $Y=1360 $dt=0
M1 7 A1 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1730 $Y=1360 $dt=0
M2 Y B0 7 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2570 $Y=1360 $dt=0
M3 8 A0 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1290 $Y=3560 $dt=1
M4 Y A1 8 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1730 $Y=3560 $dt=1
M5 VDD B0 Y VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2570 $Y=3560 $dt=1
.ends OAI21XL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AOI221XL                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AOI221XL A0 A1 VDD VSS Y B0 B1 C0
** N=12 EP=8 FDC=10
M0 9 A0 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1070 $Y=800 $dt=0
M1 Y A1 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1510 $Y=800 $dt=0
M2 10 B1 Y VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3050 $Y=800 $dt=0
M3 VSS B0 10 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3490 $Y=800 $dt=0
M4 Y C0 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=4330 $Y=800 $dt=0
M5 12 A0 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=670 $Y=3180 $dt=1
M6 VDD A1 12 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1510 $Y=3180 $dt=1
M7 12 B1 11 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3050 $Y=2840 $dt=1
M8 11 B0 12 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3890 $Y=2840 $dt=1
M9 Y C0 11 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=4730 $Y=2840 $dt=1
.ends AOI221XL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OAI222XL                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OAI222XL A1 A0 VDD VSS Y B0 C0 B1 C1
** N=14 EP=9 FDC=12
M0 10 A0 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=610 $Y=1320 $dt=0
M1 VSS A1 10 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1450 $Y=1320 $dt=0
M2 10 B1 11 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2950 $Y=1200 $dt=0
M3 11 B0 10 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3790 $Y=1200 $dt=0
M4 Y C0 11 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=4630 $Y=1200 $dt=0
M5 11 C1 Y VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=5470 $Y=1200 $dt=0
M6 12 A0 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1010 $Y=3700 $dt=1
M7 Y A1 12 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1450 $Y=3700 $dt=1
M8 13 B1 Y VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2950 $Y=3700 $dt=1
M9 VDD B0 13 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3790 $Y=3700 $dt=1
M10 14 C0 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=4630 $Y=3700 $dt=1
M11 Y C1 14 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=5070 $Y=3700 $dt=1
.ends OAI222XL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MXI2XL                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MXI2XL Y A VDD VSS S0 B
** N=11 EP=6 FDC=10
M0 8 A VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=720 $Y=1320 $dt=0
M1 Y 7 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1160 $Y=1320 $dt=0
M2 9 S0 Y VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2000 $Y=1320 $dt=0
M3 VSS B 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2460 $Y=1320 $dt=0
M4 7 S0 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3300 $Y=1320 $dt=0
M5 10 A VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=720 $Y=3700 $dt=1
M6 Y S0 10 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1160 $Y=3700 $dt=1
M7 11 7 Y VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2000 $Y=3700 $dt=1
M8 VDD B 11 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2440 $Y=3700 $dt=1
M9 7 S0 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3280 $Y=3700 $dt=1
.ends MXI2XL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: CLKXOR2X1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt CLKXOR2X1 Y VDD VSS A B
** N=10 EP=5 FDC=12
M0 VSS 8 Y VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=710 $Y=980 $dt=0
M1 6 A VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1830 $Y=1080 $dt=0
M2 8 7 6 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3110 $Y=1080 $dt=0
M3 9 B 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3950 $Y=1080 $dt=0
M4 VSS 6 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=4390 $Y=1080 $dt=0
M5 7 B VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=5230 $Y=1080 $dt=0
M6 VDD 8 Y VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=780 $Y=3120 $dt=1
M7 6 A VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1860 $Y=3240 $dt=1
M8 8 B 6 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2700 $Y=3240 $dt=1
M9 10 7 8 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3540 $Y=3240 $dt=1
M10 VDD 6 10 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=4150 $Y=3240 $dt=1
M11 7 B VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=4990 $Y=3240 $dt=1
.ends CLKXOR2X1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: TBUFX1                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt TBUFX1 OE A VDD VSS Y
** N=10 EP=5 FDC=12
M0 9 OE 6 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=720 $Y=1240 $dt=0
M1 VSS A 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1160 $Y=1240 $dt=0
M2 8 OE VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2360 $Y=1240 $dt=0
M3 7 8 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3990 $Y=1240 $dt=0
M4 VSS A 7 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=4830 $Y=1240 $dt=0
M5 Y 7 VSS VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=5790 $Y=900 $dt=0
M6 6 OE VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=710 $Y=3460 $dt=1
M7 VDD A 6 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1550 $Y=3460 $dt=1
M8 8 OE VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2630 $Y=3460 $dt=1
M9 10 8 7 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=4370 $Y=3120 $dt=1
M10 VDD A 10 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=4810 $Y=3120 $dt=1
M11 Y 6 VDD VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=6050 $Y=3120 $dt=1
.ends TBUFX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DFFTRXL                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DFFTRXL QN VDD VSS Q CK D RN
** N=20 EP=7 FDC=30
M0 VSS 14 QN VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=710 $Y=1360 $dt=0
M1 14 12 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1550 $Y=1360 $dt=0
M2 VSS 12 Q VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3170 $Y=1340 $dt=0
M3 9 CK VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=4130 $Y=1340 $dt=0
M4 VSS 13 12 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=5750 $Y=1320 $dt=0
M5 15 12 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=6710 $Y=1320 $dt=0
M6 13 9 15 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=7230 $Y=1320 $dt=0
M7 10 8 13 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=8310 $Y=1320 $dt=0
M8 VSS 11 10 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=9150 $Y=1320 $dt=0
M9 16 10 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=10070 $Y=1320 $dt=0
M10 11 8 16 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=10510 $Y=1320 $dt=0
M11 17 9 11 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=11350 $Y=1320 $dt=0
M12 VSS 9 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=13210 $Y=1320 $dt=0
M13 18 RN VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=14150 $Y=1320 $dt=0
M14 17 D 18 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=14750 $Y=1320 $dt=0
M15 VDD 14 QN VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=710 $Y=2680 $dt=1
M16 14 12 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1550 $Y=2680 $dt=1
M17 VDD 12 Q VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3170 $Y=3180 $dt=1
M18 9 CK VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=4010 $Y=3180 $dt=1
M19 VDD 13 12 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=5630 $Y=3240 $dt=1
M20 19 12 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=6710 $Y=3240 $dt=1
M21 13 8 19 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=7150 $Y=3240 $dt=1
M22 10 9 13 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=7990 $Y=3240 $dt=1
M23 VDD 11 10 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=9030 $Y=3240 $dt=1
M24 20 10 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=10110 $Y=3240 $dt=1
M25 11 9 20 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=10550 $Y=3240 $dt=1
M26 17 8 11 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=11390 $Y=3240 $dt=1
M27 VDD 9 8 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=13150 $Y=2680 $dt=1
M28 17 RN VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=13990 $Y=2680 $dt=1
M29 VDD D 17 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=14830 $Y=2680 $dt=1
.ends DFFTRXL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND2BX1                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND2BX1 B Y VDD VSS AN
** N=7 EP=5 FDC=6
M0 7 B Y VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=1120 $Y=800 $dt=0
M1 VSS 6 7 VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=1560 $Y=800 $dt=0
M2 6 AN VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2520 $Y=1180 $dt=0
M3 Y B VDD VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=840 $Y=3120 $dt=1
M4 VDD 6 Y VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=1680 $Y=3120 $dt=1
M5 6 AN VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2520 $Y=3240 $dt=1
.ends NAND2BX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DFFSHQX1                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DFFSHQX1 Q VDD VSS SN D CK
** N=20 EP=6 FDC=28
M0 VSS 11 Q VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=1280 $Y=900 $dt=0
M1 VSS 12 11 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=2900 $Y=880 $dt=0
M2 13 SN VSS VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=3740 $Y=880 $dt=0
M3 14 11 13 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=4540 $Y=880 $dt=0
M4 12 7 14 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=4980 $Y=880 $dt=0
M5 9 8 12 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=5820 $Y=880 $dt=0
M6 VSS 7 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=8520 $Y=1100 $dt=0
M7 15 SN VSS VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=9510 $Y=980 $dt=0
M8 9 10 15 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=9950 $Y=980 $dt=0
M9 16 9 VSS VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=11990 $Y=800 $dt=0
M10 10 8 16 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=12630 $Y=800 $dt=0
M11 17 7 10 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=13750 $Y=800 $dt=0
M12 VSS D 17 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=14190 $Y=800 $dt=0
M13 7 CK VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=15030 $Y=1000 $dt=0
M14 VDD 11 Q VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=1280 $Y=2680 $dt=1
M15 VDD 12 11 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=2900 $Y=3380 $dt=1
M16 18 SN VDD VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=3740 $Y=3380 $dt=1
M17 VDD 11 18 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=4580 $Y=3380 $dt=1
M18 12 8 18 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=6360 $Y=3380 $dt=1
M19 9 7 12 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=7200 $Y=3380 $dt=1
M20 VDD 7 8 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=8910 $Y=2900 $dt=1
M21 9 SN VDD VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=10110 $Y=2900 $dt=1
M22 VDD 10 9 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=10950 $Y=2900 $dt=1
M23 19 9 VDD VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=11910 $Y=2900 $dt=1
M24 10 7 19 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=12510 $Y=2900 $dt=1
M25 20 8 10 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=13350 $Y=3000 $dt=1
M26 VDD D 20 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=13790 $Y=3000 $dt=1
M27 7 CK VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=14630 $Y=3320 $dt=1
.ends DFFSHQX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: SDFFQX1                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt SDFFQX1 Q CK VDD VSS D SE SI
** N=23 EP=7 FDC=32
M0 VSS 13 Q VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=710 $Y=980 $dt=0
M1 10 CK VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1670 $Y=1360 $dt=0
M2 VSS 14 13 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3290 $Y=1360 $dt=0
M3 15 13 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=4350 $Y=1360 $dt=0
M4 14 10 15 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=5030 $Y=1360 $dt=0
M5 11 9 14 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=5870 $Y=1360 $dt=0
M6 VSS 12 11 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=7030 $Y=1360 $dt=0
M7 16 11 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=7910 $Y=1360 $dt=0
M8 12 9 16 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=8350 $Y=1360 $dt=0
M9 17 10 12 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=9190 $Y=1360 $dt=0
M10 VSS 10 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=11050 $Y=820 $dt=0
M11 18 D VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=11890 $Y=820 $dt=0
M12 17 8 18 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=12330 $Y=820 $dt=0
M13 19 SE 17 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=13170 $Y=820 $dt=0
M14 VSS SI 19 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=13610 $Y=820 $dt=0
M15 8 SE VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=14450 $Y=820 $dt=0
M16 VDD 13 Q VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=710 $Y=3120 $dt=1
M17 10 CK VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1670 $Y=3120 $dt=1
M18 VDD 14 13 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3630 $Y=3200 $dt=1
M19 20 13 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=4710 $Y=3200 $dt=1
M20 14 9 20 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=5150 $Y=3200 $dt=1
M21 11 10 14 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=5990 $Y=3200 $dt=1
M22 VDD 12 11 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=6830 $Y=3200 $dt=1
M23 21 11 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=7910 $Y=3200 $dt=1
M24 12 10 21 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=8350 $Y=3200 $dt=1
M25 17 9 12 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=9230 $Y=3200 $dt=1
M26 VDD 10 9 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=11050 $Y=3700 $dt=1
M27 22 D VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=11890 $Y=3700 $dt=1
M28 17 SE 22 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=12330 $Y=3700 $dt=1
M29 23 8 17 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=13170 $Y=3700 $dt=1
M30 VDD SI 23 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=13610 $Y=3700 $dt=1
M31 8 SE VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=14450 $Y=3700 $dt=1
.ends SDFFQX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AOI21XL                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AOI21XL A0 A1 VDD VSS B0 Y
** N=8 EP=6 FDC=6
M0 7 A0 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1130 $Y=880 $dt=0
M1 Y A1 7 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1730 $Y=880 $dt=0
M2 VSS B0 Y VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2570 $Y=880 $dt=0
M3 VDD A0 8 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=710 $Y=2920 $dt=1
M4 8 A1 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1730 $Y=2920 $dt=1
M5 Y B0 8 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2570 $Y=2920 $dt=1
.ends AOI21XL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INVXL                                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INVXL A Y VDD VSS
** N=4 EP=4 FDC=2
M0 Y A VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=710 $Y=1360 $dt=0
M1 Y A VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=710 $Y=2910 $dt=1
.ends INVXL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INVX1                                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INVX1 Y A VDD VSS
** N=4 EP=4 FDC=2
M0 Y A VSS VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=710 $Y=870 $dt=0
M1 Y A VDD VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=710 $Y=2680 $dt=1
.ends INVX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: controller1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt controller1 VDD VSS clk dataout[0] dataout[1] dataout[2] dataout[3] dataout[4] dataout[5] dataout[6]
+ dataout[7] rst status
** N=51 EP=13 FDC=256
X0 1 2 3 VDD VSS 6 NAND3BX1 $T=69600 84100 1 180 $X=64360 $Y=83740
X1 7 8 VDD VSS CLKINVX1 $T=44080 31900 0 0 $X=43480 $Y=31540
X2 dataout[5] 10 VDD VSS CLKINVX1 $T=64960 84100 1 180 $X=62620 $Y=83740
X3 11 12 VDD VSS CLKINVX1 $T=66700 84100 0 180 $X=64360 $Y=78280
X4 dataout[2] 3 VDD VSS CLKINVX1 $T=69600 84100 0 0 $X=69000 $Y=83740
X5 dataout[4] 15 16 17 VDD VSS 12 OAI211XL $T=85260 84100 0 180 $X=80600 $Y=78280
X6 dataout[7] 19 20 21 VDD VSS 1 AOI211XL $T=75400 84100 1 180 $X=70740 $Y=83740
X7 dataout[4] 22 23 15 VDD VSS 24 AOI211XL $T=82360 84100 0 0 $X=81760 $Y=83740
X8 dataout[7] 25 VDD VSS 21 24 OAI21XL $T=77720 84100 0 0 $X=77120 $Y=83740
X9 dataout[0] 12 VDD VSS 2 dataout[3] 28 29 AOI221XL $T=56840 84100 1 180 $X=50440 $Y=83740
X10 30 10 VDD VSS 6 dataout[3] 12 31 dataout[0] OAI222XL $T=63220 84100 1 180 $X=56240 $Y=83740
X11 29 32 VDD VSS dataout[1] 34 MXI2XL $T=51040 84100 1 180 $X=45800 $Y=83740
X12 22 VDD VSS dataout[6] 36 CLKXOR2X1 $T=87580 84100 1 0 $X=86980 $Y=78280
X13 37 38 VDD VSS 34 TBUFX1 $T=51040 31900 0 180 $X=43480 $Y=26080
X14 37 38 VDD VSS 39 TBUFX1 $T=49880 31900 0 0 $X=49280 $Y=31540
X15 37 38 VDD VSS 36 TBUFX1 $T=49880 42340 1 0 $X=49280 $Y=36520
X16 37 38 VDD VSS 30 TBUFX1 $T=59740 31900 0 0 $X=59140 $Y=31540
X17 37 38 VDD VSS 11 TBUFX1 $T=59740 42340 1 0 $X=59140 $Y=36520
X18 37 VDD VSS 40 clk 8 42 DFFTRXL $T=52200 31900 1 0 $X=51600 $Y=26080
X19 43 7 VDD VSS rst NAND2BX1 $T=38860 31900 1 180 $X=34780 $Y=31540
X20 43 VDD VSS 45 46 clk DFFSHQX1 $T=27260 31900 1 0 $X=26660 $Y=26080
X21 38 clk VDD VSS 38 8 47 SDFFQX1 $T=59160 21460 1 180 $X=42900 $Y=21100
X22 48 49 VDD VSS 50 46 AOI21XL $T=38280 21460 1 180 $X=34200 $Y=21100
X23 rst 45 VDD VSS INVXL $T=35380 31900 1 180 $X=33040 $Y=31540
X24 50 43 VDD VSS INVX1 $T=33060 21460 0 0 $X=32460 $Y=21100
.ends controller1
